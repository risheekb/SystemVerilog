module top;
  import uvm_pkg::*;
  import hello::*;

  initial run_test();
endmodule
