/***********************************************************************
 * Example UVM Testbench to verify an Instruction Register design.
 *
 * Class: lab_driver
 *
 * Defines a driver component within the UVM testbench.
 * Requests transactions from a sequence and drives the DUT ports
 * with those transaction values via a virtual interface to the DUT.
 ***********************************************************************
 * Copyright 2016-2023 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 *
 * CBS 191212 - Switched to drv_bfm
 * CBS 170714 - Cleaned up
 **********************************************************************/

`ifndef lab_driver_exists
 `define lab_driver_exists


class lab_driver extends uvm_driver #(lab_tx_in);

  // Register this class name in the factory
  `uvm_component_utils(lab_driver)
  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  lab_tx_agent_config tx_cfg;
  virtual tx_driver_bfm drv_bfm;   // virtual interface pointer

  virtual function void build_phase(uvm_phase phase);
    // Fetch the agent configuration
    // You will learn about the uvm_config_db in Lab 8
    if (!uvm_config_db #(lab_tx_agent_config)::get(this, "", "tx_cfg", tx_cfg))
      `uvm_fatal(get_type_name(), "Failed to get tx_cfg from uvm_config_db")
    drv_bfm = tx_cfg.drv_bfm;
  endfunction: build_phase


  //
  // LAB 4 ASSIGNMENT:
  // Add the run_phase() task that:
  // 1) Declares a lab_tx_in sequence_item handle
  // 2) Contains a forever loop that:
  //    - Calls get_next_item(tx) to request a sequence_item object.
  //    - Calls a drv_bfm.send(tx) task to drive the sequence_item values
  //    - Calls item_done() to release the sequence item
  //
  //ADD YOUR CODE HERE...
  //BEGIN SOLUTION
  virtual task run_phase(uvm_phase phase);
    forever begin
      lab_tx_in tx;

      seq_item_port.get_next_item(tx);
      drv_bfm.send(.reset_n(tx.reset_n),
		   .load_en(tx.load_en),
		   .read_pointer(tx.read_pointer),
		   .write_pointer(tx.write_pointer),
		   .operand_a(tx.operand_a),
		   .operand_b(tx.operand_b),
		   .opcode(tx.opcode));
      seq_item_port.item_done();
    end
  endtask: run_phase
  //END SOLUTION



endclass: lab_driver
`endif
