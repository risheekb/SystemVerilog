/***********************************************************************
 * Example to show compare() and do_compare() functions
 * Compile & run with compile script or:
 * % qrun tx_pkg.sv seq_item.sv
 ***********************************************************************
 * Copyright 2016-2023 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/

module seq_item;
  timeunit 1ns/1ns;
`include "uvm_macros.svh"
  import uvm_pkg::*;
  import tx_pkg::*;

  initial begin
    $timeformat(-9, 0, "ns", 0);
    run_test("seq_item_test");
  end

endmodule : seq_item
