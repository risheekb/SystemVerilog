package ram_pkg;
  parameter DEPTH = 16;
  parameter ADDR_WIDTH = $clog2(DEPTH);
  parameter DATA_WIDTH = 16;
endpackage
