class apb_cov;
  task run();
    $display("apb_cov::run");
  endtask
endclass
