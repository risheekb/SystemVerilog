/***********************************************************************
 * Transaction for TX UVM example
 ***********************************************************************
 * Copyright 2016-2023 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/

class tx_item extends uvm_sequence_item;
  `uvm_object_utils(tx_item);
  function new(string name="tx_item");
    super.new(name);
  endfunction : new

  rand bit [7:0] data;

endclass

typedef uvm_sequencer #(tx_item) tx_sequencer;
