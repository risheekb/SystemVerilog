package noise_pkg;
  import uvm_pkg::*;
`include "uvm_macros.svh"

`include "agt_config.svh"

`include "main_sequence.svh"
`include "noise_sequence.svh"
`include "two_vseq.svh"

`include "multi_agt.svh"
`include "multi_env.svh"
`include "multi_test.svh"
endpackage : noise_pkg
