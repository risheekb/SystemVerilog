class apb_mon;
  task run();
    $display("apb_mon::run");
  endtask
endclass

