class axi_responder;
  task run();
    $display("axi_responder::run");
  endtask
endclass
