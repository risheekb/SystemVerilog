class dma_ref;
  task run();
    $display("dma_ref::run");
  endtask
endclass
