/***********************************************************************
 * HVL top for UVM configuration flow example
 ***********************************************************************
 * Copyright 2016-2017 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/

module top_tb;
   import uvm_pkg::*;
   import spi_pkg::*;
   import usb_pkg::*;

   initial begin
//      $timeformat(-9,0,"ns",3); // Shorten messages on slides
      run_test();
   end

  initial #1000ns $fatal(0, "Time out!");

endmodule
