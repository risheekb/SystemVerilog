interface axi_inf(input clk,reset);

  bit [`ID_BITS-1:0]               AWID0;
  bit [32-1:0]                     AWADDR0;
  bit [`LEN_BITS-1:0]              AWLEN0;
  bit [`SIZE_BITS-1:0]             AWSIZE0;
  bit                              AWVALID0;
  bit                              AWREADY0;
  bit [`ID_BITS-1:0]               WID0;
  bit [64-1:0]                     WDATA0;
  bit [64/8-1:0]                   WSTRB0;
  bit                              WLAST0;
  bit                              WVALID0;
  bit                              WREADY0;
  bit [`ID_BITS-1:0]               BID0;
  bit [1:0]                        BRESP0;
  bit                              BVALID0;
  bit                              BREADY0;
  bit [`ID_BITS-1:0]               ARID0;
  bit [32-1:0]                     ARADDR0;
  bit [`LEN_BITS-1:0]              ARLEN0;
  bit [`SIZE_BITS-1:0]             ARSIZE0;
  bit                              ARVALID0;
  bit                              ARREADY0;
  bit [`ID_BITS-1:0]               RID0;
  bit [64-1:0]                     RDATA0;
  bit [1:0]                        RRESP0;
  bit                              RLAST0;
  bit                              RVALID0;
  bit                              RREADY0;

  clocking slave_cb @(posedge clk);
    default input #0;
    default output #1;
    output                         AWID0;
    output                         AWADDR0;
    output                         AWLEN0;
    output                         AWSIZE0;
    output                         AWVALID0;
    input                          AWREADY0;
    output                         WID0;
    output                         WDATA0;
    output                         WSTRB0;
    output                         WLAST0;
    output                         WVALID0;
    input                          WREADY0;
    input                          BID0;
    input                          BRESP0;
    input                          BVALID0;
    output                         BREADY0;
    output                         ARID0;
    output                         ARADDR0;
    output                         ARLEN0;
    output                         ARSIZE0;
    output                         ARVALID0;
    input                          ARREADY0;
    input                          RID0;
    input                          RDATA0;
    input                          RRESP0;
    input                          RLAST0;
    input                          RVALID0;
    output                         RREADY0;
  endclocking

  clocking monitor_cb @(posedge clk);
    default input #0;
    input                         AWID0;
    input                         AWADDR0;
    input                         AWLEN0;
    input                         AWSIZE0;
    input                         AWVALID0;
    input                          AWREADY0;
    input                         WID0;
    input                         WDATA0;
    input                         WSTRB0;
    input                         WLAST0;
    input                         WVALID0;
    input                          WREADY0;
    input                          BID0;
    input                          BRESP0;
    input                          BVALID0;
    input                         BREADY0;
    input                         ARID0;
    input                         ARADDR0;
    input                         ARLEN0;
    input                         ARSIZE0;
    input                         ARVALID0;
    input                          ARREADY0;
    input                          RID0;
    input                          RDATA0;
    input                          RRESP0;
    input                          RLAST0;
    input                          RVALID0;
    input                         RREADY0;
  endclocking

  modport slave_mp(clocking slave_cb);
  modport monitor_mp(clocking monitor_mp);
endinterface
