class apb_cov;
  apb_tx tx_h;
  covergroup apb_cg;

    CP_ADDR:coverpoint tx_h.addr{

      //CH0 REGISTERS//
      bins CH0_CMD_REG0            ={`CH0_CMD_REG0};
      bins CH0_CMD_REG1            ={`CH0_CMD_REG1};
      bins CH0_CMD_REG2            ={`CH0_CMD_REG2};
      bins CH0_CMD_REG3            ={`CH0_CMD_REG3};
      bins CH0_STATIC_REG0         ={`CH0_STATIC_REG0};
      bins CH0_STATIC_REG1         ={`CH0_STATIC_REG1};
      bins CH0_STATIC_REG2         ={`CH0_STATIC_REG2};
      bins CH0_STATIC_REG3         ={`CH0_STATIC_REG3};
      bins CH0_STATIC_REG4         ={`CH0_STATIC_REG4};
      bins CH0_RESTRICT_REG        ={`CH0_RESTRICT_REG};
      bins CH0_READ_OFFSET_REG     ={`CH0_READ_OFFSET_REG};
      bins CH0_WRITE_OFFSET_REG    ={`CH0_WRITE_OFFSET_REG};
      bins CH0_FIFO_FULLNESS_REG   ={`CH0_FIFO_FULLNESS_REG};
      bins CH0_CMD_OUTS_REG            ={`CH0_CMD_OUTS_REG};
      bins CH0_CH_ENABLE_REG       ={`CH0_CH_ENABLE_REG};
      bins CH0_CH_START_REG        ={`CH0_CH_START_REG};
      bins CH0_CH_ACTIVE_REG       ={`CH0_CH_ACTIVE_REG};
      bins CH0_COUNT_REG           ={`CH0_COUNT_REG};
      bins CH0_INT_RAWSTAT_REG     ={`CH0_INT_RAWSTAT_REG};
      bins CH0_INT_CLEAR_REG       ={`CH0_INT_CLEAR_REG};
      bins CH0_INT_ENABLE_REG      ={`CH0_INT_ENABLE_REG};
      bins CH0_INT_STATUS_REG      ={`CH0_INT_STATUS_REG};
      //CHANNEL 1 REGISTERS
      bins CH1_CMD_REG0            ={`CH1_CMD_REG0};
      bins CH1_CMD_REG1            ={`CH1_CMD_REG1};
      bins CH1_CMD_REG2            ={`CH1_CMD_REG2};
      bins CH1_CMD_REG3            ={`CH1_CMD_REG3};
      bins CH1_STATIC_REG0         ={`CH1_STATIC_REG0};
      bins CH1_STATIC_REG1         ={`CH1_STATIC_REG1};
      bins CH1_STATIC_REG2         ={`CH1_STATIC_REG2};
      bins CH1_STATIC_REG3         ={`CH1_STATIC_REG3};
      bins CH1_STATIC_REG4         ={`CH1_STATIC_REG4};
      bins CH1_RESTRICT_REG        ={`CH1_RESTRICT_REG};
      bins CH1_READ_OFFSET_REG     ={`CH1_READ_OFFSET_REG};
      bins CH1_WRITE_OFFSET_REG    ={`CH1_WRITE_OFFSET_REG};
      bins CH1_FIFO_FULLNESS_REG   ={`CH1_FIFO_FULLNESS_REG};
      bins CH1_CMD_OUTS_REG            ={`CH1_CMD_OUTS_REG};
      bins CH1_CH_ENABLE_REG       ={`CH1_CH_ENABLE_REG};
      bins CH1_CH_START_REG        ={`CH1_CH_START_REG};
      bins CH1_CH_ACTIVE_REG       ={`CH1_CH_ACTIVE_REG};
      bins CH1_COUNT_REG           ={`CH1_COUNT_REG};
      bins CH1_INT_RAWSTAT_REG     ={`CH1_INT_RAWSTAT_REG};
      bins CH1_INT_CLEAR_REG       ={`CH1_INT_CLEAR_REG};
      bins CH1_INT_ENABLE_REG      ={`CH1_INT_ENABLE_REG};
      bins CH1_INT_STATUS_REG      ={`CH1_INT_STATUS_REG};
      //CHANNEL 2 REGISTERS
      bins CH2_CMD_REG0            ={`CH2_CMD_REG0};
      bins CH2_CMD_REG1            ={`CH2_CMD_REG1};
      bins CH2_CMD_REG2            ={`CH2_CMD_REG2};
      bins CH2_CMD_REG3            ={`CH2_CMD_REG3};
      bins CH2_STATIC_REG0         ={`CH2_STATIC_REG0};
      bins CH2_STATIC_REG1         ={`CH2_STATIC_REG1};
      bins CH2_STATIC_REG2         ={`CH2_STATIC_REG2};
      bins CH2_STATIC_REG3         ={`CH2_STATIC_REG3};
      bins CH2_STATIC_REG4         ={`CH2_STATIC_REG4};
      bins CH2_RESTRICT_REG        ={`CH2_RESTRICT_REG};
      bins CH2_READ_OFFSET_REG     ={`CH2_READ_OFFSET_REG};
      bins CH2_WRITE_OFFSET_REG    ={`CH2_WRITE_OFFSET_REG};
      bins CH2_FIFO_FULLNESS_REG   ={`CH2_FIFO_FULLNESS_REG};
      bins CH2_CMD_OUTS_REG            ={`CH2_CMD_OUTS_REG};
      bins CH2_CH_ENABLE_REG       ={`CH2_CH_ENABLE_REG};
      bins CH2_CH_START_REG        ={`CH2_CH_START_REG};
      bins CH2_CH_ACTIVE_REG       ={`CH2_CH_ACTIVE_REG};
      bins CH2_COUNT_REG           ={`CH2_COUNT_REG};
      bins CH2_INT_RAWSTAT_REG     ={`CH2_INT_RAWSTAT_REG};
      bins CH2_INT_CLEAR_REG       ={`CH2_INT_CLEAR_REG};
      bins CH2_INT_ENABLE_REG      ={`CH2_INT_ENABLE_REG};
      bins CH2_INT_STATUS_REG      ={`CH2_INT_STATUS_REG};
      //CHANNEL 3 REGISTERS
      bins CH3_CMD_REG0            ={`CH3_CMD_REG0};
      bins CH3_CMD_REG1            ={`CH3_CMD_REG1};
      bins CH3_CMD_REG2            ={`CH3_CMD_REG2};
      bins CH3_CMD_REG3            ={`CH3_CMD_REG3};
      bins CH3_STATIC_REG0         ={`CH3_STATIC_REG0};
      bins CH3_STATIC_REG1         ={`CH3_STATIC_REG1};
      bins CH3_STATIC_REG2         ={`CH3_STATIC_REG2};
      bins CH3_STATIC_REG3         ={`CH3_STATIC_REG3};
      bins CH3_STATIC_REG4         ={`CH3_STATIC_REG4};
      bins CH3_RESTRICT_REG        ={`CH3_RESTRICT_REG};
      bins CH3_READ_OFFSET_REG     ={`CH3_READ_OFFSET_REG};
      bins CH3_WRITE_OFFSET_REG    ={`CH3_WRITE_OFFSET_REG};
      bins CH3_FIFO_FULLNESS_REG   ={`CH3_FIFO_FULLNESS_REG};
      bins CH3_CMD_OUTS_REG            ={`CH3_CMD_OUTS_REG};
      bins CH3_CH_ENABLE_REG       ={`CH3_CH_ENABLE_REG};
      bins CH3_CH_START_REG        ={`CH3_CH_START_REG};
      bins CH3_CH_ACTIVE_REG       ={`CH3_CH_ACTIVE_REG};
      bins CH3_COUNT_REG           ={`CH3_COUNT_REG};
      bins CH3_INT_RAWSTAT_REG     ={`CH3_INT_RAWSTAT_REG};
      bins CH3_INT_CLEAR_REG       ={`CH3_INT_CLEAR_REG};
      bins CH3_INT_ENABLE_REG      ={`CH3_INT_ENABLE_REG};
      bins CH3_INT_STATUS_REG      ={`CH3_INT_STATUS_REG};
      //CHANNEL 4 REGISTERS
      bins CH4_CMD_REG0            ={`CH4_CMD_REG0};
      bins CH4_CMD_REG1            ={`CH4_CMD_REG1};
      bins CH4_CMD_REG2            ={`CH4_CMD_REG2};
      bins CH4_CMD_REG3            ={`CH4_CMD_REG3};
      bins CH4_STATIC_REG0         ={`CH4_STATIC_REG0};
      bins CH4_STATIC_REG1         ={`CH4_STATIC_REG1};
      bins CH4_STATIC_REG2         ={`CH4_STATIC_REG2};
      bins CH4_STATIC_REG3         ={`CH4_STATIC_REG3};
      bins CH4_STATIC_REG4         ={`CH4_STATIC_REG4};
      bins CH4_RESTRICT_REG        ={`CH4_RESTRICT_REG};
      bins CH4_READ_OFFSET_REG     ={`CH4_READ_OFFSET_REG};
      bins CH4_WRITE_OFFSET_REG    ={`CH4_WRITE_OFFSET_REG};
      bins CH4_FIFO_FULLNESS_REG   ={`CH4_FIFO_FULLNESS_REG};
      bins CH4_CMD_OUTS_REG            ={`CH4_CMD_OUTS_REG};
      bins CH4_CH_ENABLE_REG       ={`CH4_CH_ENABLE_REG};
      bins CH4_CH_START_REG        ={`CH4_CH_START_REG};
      bins CH4_CH_ACTIVE_REG       ={`CH4_CH_ACTIVE_REG};
      bins CH4_COUNT_REG           ={`CH4_COUNT_REG};
      bins CH4_INT_RAWSTAT_REG     ={`CH4_INT_RAWSTAT_REG};
      bins CH4_INT_CLEAR_REG       ={`CH4_INT_CLEAR_REG};
      bins CH4_INT_ENABLE_REG      ={`CH4_INT_ENABLE_REG};
      bins CH4_INT_STATUS_REG      ={`CH4_INT_STATUS_REG};
      //CHANNEL 5 REGISTERS
      bins CH5_CMD_REG0            ={`CH5_CMD_REG0};
      bins CH5_CMD_REG1            ={`CH5_CMD_REG1};
      bins CH5_CMD_REG2            ={`CH5_CMD_REG2};
      bins CH5_CMD_REG3            ={`CH5_CMD_REG3};
      bins CH5_STATIC_REG0         ={`CH5_STATIC_REG0};
      bins CH5_STATIC_REG1         ={`CH5_STATIC_REG1};
      bins CH5_STATIC_REG2         ={`CH5_STATIC_REG2};
      bins CH5_STATIC_REG3         ={`CH5_STATIC_REG3};
      bins CH5_STATIC_REG4         ={`CH5_STATIC_REG4};
      bins CH5_RESTRICT_REG        ={`CH5_RESTRICT_REG};
      bins CH5_READ_OFFSET_REG     ={`CH5_READ_OFFSET_REG};
      bins CH5_WRITE_OFFSET_REG    ={`CH5_WRITE_OFFSET_REG};
      bins CH5_FIFO_FULLNESS_REG   ={`CH5_FIFO_FULLNESS_REG};
      bins CH5_CMD_OUTS_REG            ={`CH5_CMD_OUTS_REG};
      bins CH5_CH_ENABLE_REG       ={`CH5_CH_ENABLE_REG};
      bins CH5_CH_START_REG        ={`CH5_CH_START_REG};
      bins CH5_CH_ACTIVE_REG       ={`CH5_CH_ACTIVE_REG};
      bins CH5_COUNT_REG           ={`CH5_COUNT_REG};
      bins CH5_INT_RAWSTAT_REG     ={`CH5_INT_RAWSTAT_REG};
      bins CH5_INT_CLEAR_REG       ={`CH5_INT_CLEAR_REG};
      bins CH5_INT_ENABLE_REG      ={`CH5_INT_ENABLE_REG};
      bins CH5_INT_STATUS_REG      ={`CH5_INT_STATUS_REG};
      //CHANNEL 6 REGISTERS
      bins CH6_CMD_REG0            ={`CH6_CMD_REG0};
      bins CH6_CMD_REG1            ={`CH6_CMD_REG1};
      bins CH6_CMD_REG2            ={`CH6_CMD_REG2};
      bins CH6_CMD_REG3            ={`CH6_CMD_REG3};
      bins CH6_STATIC_REG0         ={`CH6_STATIC_REG0};
      bins CH6_STATIC_REG1         ={`CH6_STATIC_REG1};
      bins CH6_STATIC_REG2         ={`CH6_STATIC_REG2};
      bins CH6_STATIC_REG3         ={`CH6_STATIC_REG3};
      bins CH6_STATIC_REG4         ={`CH6_STATIC_REG4};
      bins CH6_RESTRICT_REG        ={`CH6_RESTRICT_REG};
      bins CH6_READ_OFFSET_REG     ={`CH6_READ_OFFSET_REG};
      bins CH6_WRITE_OFFSET_REG    ={`CH6_WRITE_OFFSET_REG};
      bins CH6_FIFO_FULLNESS_REG   ={`CH6_FIFO_FULLNESS_REG};
      bins CH6_CMD_OUTS_REG            ={`CH6_CMD_OUTS_REG};
      bins CH6_CH_ENABLE_REG       ={`CH6_CH_ENABLE_REG};
      bins CH6_CH_START_REG        ={`CH6_CH_START_REG};
      bins CH6_CH_ACTIVE_REG       ={`CH6_CH_ACTIVE_REG};
      bins CH6_COUNT_REG           ={`CH6_COUNT_REG};
      bins CH6_INT_RAWSTAT_REG     ={`CH6_INT_RAWSTAT_REG};
      bins CH6_INT_CLEAR_REG       ={`CH6_INT_CLEAR_REG};
      bins CH6_INT_ENABLE_REG      ={`CH6_INT_ENABLE_REG};
      bins CH6_INT_STATUS_REG      ={`CH6_INT_STATUS_REG};
      //CHANNEL 7 REGISTERS
      bins CH7_CMD_REG0            ={`CH7_CMD_REG0};
      bins CH7_CMD_REG1            ={`CH7_CMD_REG1};
      bins CH7_CMD_REG2            ={`CH7_CMD_REG2};
      bins CH7_CMD_REG3            ={`CH7_CMD_REG3};
      bins CH7_STATIC_REG0         ={`CH7_STATIC_REG0};
      bins CH7_STATIC_REG1         ={`CH7_STATIC_REG1};
      bins CH7_STATIC_REG2         ={`CH7_STATIC_REG2};
      bins CH7_STATIC_REG3         ={`CH7_STATIC_REG3};
      bins CH7_STATIC_REG4         ={`CH7_STATIC_REG4};
      bins CH7_RESTRICT_REG        ={`CH7_RESTRICT_REG};
      bins CH7_READ_OFFSET_REG     ={`CH7_READ_OFFSET_REG};
      bins CH7_WRITE_OFFSET_REG    ={`CH7_WRITE_OFFSET_REG};
      bins CH7_FIFO_FULLNESS_REG   ={`CH7_FIFO_FULLNESS_REG};
      bins CH7_CMD_OUTS_REG            ={`CH7_CMD_OUTS_REG};
      bins CH7_CH_ENABLE_REG       ={`CH7_CH_ENABLE_REG};
      bins CH7_CH_START_REG        ={`CH7_CH_START_REG};
      bins CH7_CH_ACTIVE_REG       ={`CH7_CH_ACTIVE_REG};
      bins CH7_COUNT_REG           ={`CH7_COUNT_REG};
      bins CH7_INT_RAWSTAT_REG     ={`CH7_INT_RAWSTAT_REG};
      bins CH7_INT_CLEAR_REG       ={`CH7_INT_CLEAR_REG};
      bins CH7_INT_ENABLE_REG      ={`CH7_INT_ENABLE_REG};
      bins CH7_INT_STATUS_REG      ={`CH7_INT_STATUS_REG};
      //SHARED REGISTERS
      bins INT0_STATUS             ={`INT0_STATUS};
      bins INT1_STATUS             ={`INT1_STATUS};
      bins INT2_STATUS             ={`INT2_STATUS};
      bins INT3_STATUS             ={`INT3_STATUS};
      bins INT4_STATUS             ={`INT4_STATUS};
      bins INT5_STATUS             ={`INT5_STATUS};
      bins INT6_STATUS             ={`INT6_STATUS};
      bins INT7_STATUS             ={`INT7_STATUS};
      bins CORE0_JOINT_MODE        ={`CORE0_JOINT_MODE};
      bins CORE1_JOINT_MODE        ={`CORE1_JOINT_MODE};
      bins CORE0_PRIORITY          ={`CORE0_PRIORITY};
      bins CORE1_PRIORITY          ={`CORE1_PRIORITY};
      bins CORE0_CLKDIV            ={`CORE0_CLKDIV};
      bins CORE1_CLKDIV            ={`CORE1_CLKDIV};
      bins CORE0_CH_START          ={`CORE0_CH_START};
      bins PERIPH_RX_CTRL          ={`PERIPH_RX_CTRL};
      bins PERIPH_TX_CTRL          ={`PERIPH_TX_CTRL};
      bins IDLE                    ={`IDLE};
      bins USER_DEF_STATUS         ={`USER_DEF_STATUS};
      bins USER_CORE0_DEF_STATUS0  ={`USER_CORE0_DEF_STATUS0};
      bins USER_CORE0_DEF_STATUS1  ={`USER_CORE0_DEF_STATUS1};
    }
    CP_WR_RD:coverpoint tx_h.wr_rd{
      bins WR = {1'b1};
      bins RD = {1'b0};
    }
    cross CP_ADDR,CP_WR_RD;
  endgroup
  function new();
    apb_cg= new();
  endfunction
  task run();
    $display("apb_cov::run");
    forever begin
      tx_h = new();
      dma_common::mon2cov.get(tx_h);
      apb_cg.sample();
    end
  endtask
endclass

