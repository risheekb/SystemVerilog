package tx_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  typedef class tx_agent_config;
  typedef class tx_env_config;

  `include "tx_item.svh"
  `include "tx_sequence.svh"
  `include "tx_monitor.svh"
  `include "tx_driver.svh"
  `include "tx_agent_config.svh"
  `include "tx_agent.svh"
  `include "tx_env_config.svh"
  `include "tx_env.svh"
  `include "tx_test.svh"

  
endpackage
