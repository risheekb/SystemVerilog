class apb_gen;
  task run();
    $display("apb_gen::run");
  endtask
endclass
