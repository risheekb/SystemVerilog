class axi_mon;
  task run();
    $display("axi_mon::run");
  endtask
endclass
