/***********************************************************************
 * Testbench top for "dual-top" example
 * Compile with compile_dual.bat or compile_dual.do
 ***********************************************************************
 * Copyright 2016-2023 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/

module top_tb();
  timeunit 1ns/1ns;
  import uvm_pkg::*;

  initial begin
    $timeformat(-9,0,"ns",6);
    run_test();
  end

endmodule
