class dma_ckr;
  task run();
    $display("dma_ckr::run");
  endtask
endclass
