class dma_common;
  static virtual apb_inf apb_vif;
  static virtual axi_inf axi_vif;
  static virtual periph_inf periph_vif;
endclass
