/***********************************************************************
 * Package for UVM configuration flow example
 ***********************************************************************
 * Copyright 2016-2017 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/

package usb_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"

   import spi_pkg::*;

   typedef class usb_config;

   `include "usb_item.svh"
   `include "usb_sequence.svh"
   `include "usb_fixed_addr_sequence.svh"
   `include "usb_fixed_addr2_sequence.svh"
   `include "usb_config.svh"
   `include "usb_monitor.svh"
   `include "usb_driver.svh"
   `include "usb_agent.svh"
   `include "usb_cov_collect.svh"
   `include "usb_env_config.svh"
   `include "usb_env.svh"
   `include "usb_test.svh"
   `include "usb_fixed_addr_test.svh"
   `include "usb_fixed_addr2_test.svh"

endpackage : usb_pkg
