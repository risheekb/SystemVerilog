/***********************************************************************
 * HDL top of the Design Under Test
 ***********************************************************************
 * Copyright 2016-2017 Siemens
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License"); 
 * you may not use this file except in compliance with the License.  
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/


module top_hdl();
  timeunit 1ns; timeprecision 1ns;

   import alu_pkg::*;

   alu_ifc alu_if();
   alu a1(.result  (alu_if.result),
	  .a       (alu_if.a),
	  .b       (alu_if.b),
	  .opcode  (alu_if.opcode),
	  .addr_in (alu_if.addr_in),
	  .addr_out(alu_if.addr_out),
	  .clk     (alu_if.clk),
	  .reset_n (alu_if.reset_n));

endmodule : top_hdl
