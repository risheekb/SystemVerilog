class axi_cov;
  virtual task run();
    $display("axi_cov::run");
  endtask
endclass
