class apb_bfm;
  task run();
    $display("apb_bfm::run");
  endtask
endclass
